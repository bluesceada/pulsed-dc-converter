*SRC=BZT52C5V6LP;DI_BZT52C5V6LP;Diodes;Zener <=10V; 5.60V  0.250W   Diodes Inc. QFN Zener
*SYM=HZEN
.SUBCKT DI_BZT52C5V6LP  1 2
*        Terminals    A   K
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 3.31
.MODEL DF D ( IS=18.4p RS=32.7 N=1.10
+ CJO=106p VJ=0.750 M=0.330 TT=50.1n )
.MODEL DR D ( IS=3.68f RS=24.5 N=3.00 )
.ENDS
